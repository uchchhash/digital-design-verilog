`timescale 1ns/1ps

// Module: rca_3op_16bit
// Description: This module implements a 16-bit 3-operand Ripple Carry Adder (RCA).
//              It sums three 16-bit unsigned operands (A, B, C) and an initial carry-in (Cin).
//              The maximum possible sum of three 16-bit numbers plus Cin requires 18 bits.
//              This design achieves the 3-operand addition by cascading two instances of
//              the 'rca_2op_16bit' (2-operand, 16-bit) module.
//
// Inputs:
//   A    : logic [15:0] - The first 16-bit unsigned operand.
//   B    : logic [15:0] - The second 16-bit unsigned operand.
//   C    : logic [15:0] - The third 16-bit unsigned operand.
//   Cin  : logic        - The initial carry-in to the least significant bit (bit 0) of the overall addition.
//
// Outputs:
//   S    : logic [17:0] - The 18-bit result of the addition (A + B + C + Cin).
//                        S[15:0] represents the 16-bit sum.
//                        S[16] and S[17] represent the higher-order bits due to carries
//                        propagating beyond the initial 16-bit range.
//

module rca_3op_16bit (
    input  logic [15:0] A,
    input  logic [15:0] B,
    input  logic [15:0] C,
    input  logic        Cin,
    output logic [17:0] S // 18-bit output for full sum (16-bit sum + 2 bits for potential carries)
);

    // Intermediate Wire: sum_AB_intermediate
    // This wire stores the 17-bit result of the first addition: (A + B + Cin).
    // sum_AB_intermediate[15:0] holds the 16-bit sum part.
    // sum_AB_intermediate[16] holds the carry-out from bit 15, which is essentially a value at bit position 16.
    logic [16:0] sum_AB_intermediate;

    // Instance 1: RCA0 (First Stage Addition)
    // This 'rca_2op_16bit' calculates the sum of A, B, and the module's initial Cin.
    rca_2op_16bit RCA0 (
        .A   (A),                           // First 16-bit operand for this stage
        .B   (B),                           // Second 16-bit operand for this stage
        .Cin (Cin),                         // Initial carry-in for the entire 3-operand addition
        .S   (sum_AB_intermediate)          // Output of this stage (17 bits)
    );

    // Intermediate Wire: sum_ABC_lower_intermediate
    // This wire stores the 17-bit result of the second addition:
    // (sum_AB_intermediate[15:0] + C + 0 as Cin).
    // sum_ABC_lower_intermediate[15:0] holds the 16-bit sum part.
    // sum_ABC_lower_intermediate[16] holds the carry-out from bit 15 of this second addition.
    logic [16:0] sum_ABC_lower_intermediate;

    // Instance 2: RCA1 (Second Stage Addition for Lower Bits)
    // This 'rca_2op_16bit' adds the lower 16 bits of the result from RCA0
    // with the third operand C.
    // IMPORTANT: Its Cin is set to 0. The carry from RCA0 (sum_AB_intermediate[16])
    // is treated as a separate bit to be summed at position 16, not as a ripple carry-in
    // to the least significant bit (bit 0) of this RCA1.
    rca_2op_16bit RCA1 (
        .A   (sum_AB_intermediate[15:0]), // The lower 16 bits of the sum from RCA0
        .B   (C),                         // The third 16-bit operand (C)
        .Cin (1'b0),                      // Initial carry-in for this 16-bit adder is 0
        .S   (sum_ABC_lower_intermediate) // Output of this stage (17 bits)
    );

    // Final Sum Assignment: Lower 16 bits (S[15:0])
    // The lower 16 bits of the final sum are simply the sum bits from the second RCA (RCA1).
    assign S[15:0] = sum_ABC_lower_intermediate[15:0];

    // Final Sum Assignment: Higher Bits (S[16] and S[17])
    // At bit position 16, there are two potential contributions:
    // 1. `sum_AB_intermediate[16]`: The carry that was generated by RCA0 (from A+B+Cin).
    // 2. `sum_ABC_lower_intermediate[16]`: The carry that was generated by RCA1
    //    (from sum_AB_intermediate[15:0] + C).
    // These two bits effectively represent values at the $2^{16}$ position.
    // We add them together using logical operations which mimic a half-adder:
    // - The XOR operation gives the sum bit for S[16].
    // - The AND operation gives the carry-out from S[16] to S[17].

    assign S[16] = sum_AB_intermediate[16] ^ sum_ABC_lower_intermediate[16]; // Sum bit for position 16
    assign S[17] = sum_AB_intermediate[16] & sum_ABC_lower_intermediate[16]; // Carry bit to position 17

endmodule

